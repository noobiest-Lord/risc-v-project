
module half_adder(A,B,S,C);
    input A, B;
    
    output S, C;

    // declaring interim wires

    // Module initiation

    // Logic design
    // Data flow modelling
    // assign keyword
    // AND = &
    // OR = |
    // XOR = ^
    // Not = ~ 

    assign C = A & B; // basically boiling down the function to one sentence
    assign S = A ~ B;
endmodule